module MLP #(parameter N, parameter M) (


); 



endmodule