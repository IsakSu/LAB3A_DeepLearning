


module MLP(); 



endmodule